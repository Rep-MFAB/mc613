library ieee;
use ieee.std_logic_1164.all;

entity linear_regression is
	port (
		
	)
end linear_regression;

architecture behavioral of linear_regression is
begin
	
end behavioral;
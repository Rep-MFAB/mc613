library ieee;
use ieee.std_logic_1164.all;

entity loss is
	port (
		
	)
end loss;

architecture behavioral of loss is
begin
	
end loss;